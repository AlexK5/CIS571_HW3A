`timescale 1ns / 1ns

// registers are 32 bits in RV32
`define REG_SIZE 31:0

// RV opcodes are 7 bits
`define OPCODE_SIZE 6:0

`include "../hw2a/divider_unsigned.sv"
`include "../hw2b/cla.sv"

module RegFile (
    input logic [4:0] rd,
    input logic [`REG_SIZE] rd_data,
    input logic [4:0] rs1,
    output logic [`REG_SIZE] rs1_data,
    input logic [4:0] rs2,
    output logic [`REG_SIZE] rs2_data,

    input logic clk,
    input logic we,
    input logic rst
);
  localparam int NumRegs = 32;
  logic [`REG_SIZE] regs[NumRegs];
  assign regs[0] = 32'd0; // x0 is always zero
  assign rs1_data = regs[rs1]; // 1st read port
  assign rs2_data = regs[rs2]; // 2nd read port

  
  always_ff @(posedge clk) begin
    for (int i = 1; i < NumRegs; i = i + 1) begin
      if (rst) begin
        regs[i] <= 32'd0;
      end else begin
        if (we && rd == i[4:0]) begin
          regs[i] <= rd_data;
        end
      end
    end
  end
  
  
  // TODO: your code here

endmodule

module DatapathSingleCycle (
    input wire clk,
    input wire rst,
    output logic halt,
    output logic [`REG_SIZE] pc_to_imem,
    input wire [`REG_SIZE] insn_from_imem,
    // addr_to_dmem is a read-write port
    output wire [`REG_SIZE] addr_to_dmem,
    input logic [`REG_SIZE] load_data_from_dmem,
    output wire [`REG_SIZE] store_data_to_dmem,
    output wire [3:0] store_we_to_dmem
);

  // components of the instruction
  wire [6:0] insn_funct7;
  wire [4:0] insn_rs2;
  wire [4:0] insn_rs1;
  wire [2:0] insn_funct3;
  wire [4:0] insn_rd;
  wire [`OPCODE_SIZE] insn_opcode;

  // split R-type instruction - see section 2.2 of RiscV spec
  assign {insn_funct7, insn_rs2, insn_rs1, insn_funct3, insn_rd, insn_opcode} = insn_from_imem;

  // setup for I, S, B & J type instructions
  // I - short immediates and loads
  wire [11:0] imm_i;
  assign imm_i = insn_from_imem[31:20];
  wire [ 4:0] imm_shamt = insn_from_imem[24:20];

  // S - stores
  wire [11:0] imm_s;
  assign imm_s[11:5] = insn_funct7, imm_s[4:0] = insn_rd;

  // B - conditionals
  wire [12:0] imm_b;
  assign {imm_b[12], imm_b[10:5]} = insn_funct7, {imm_b[4:1], imm_b[11]} = insn_rd, imm_b[0] = 1'b0;

  // J - unconditional jumps
  wire [20:0] imm_j;
  assign {imm_j[20], imm_j[10:1], imm_j[11], imm_j[19:12], imm_j[0]} = {insn_from_imem[31:12], 1'b0};

  wire [`REG_SIZE] imm_i_sext = {{20{imm_i[11]}}, imm_i[11:0]};
  wire [`REG_SIZE] imm_s_sext = {{20{imm_s[11]}}, imm_s[11:0]};
  wire [`REG_SIZE] imm_b_sext = {{19{imm_b[12]}}, imm_b[12:0]};
  wire [`REG_SIZE] imm_j_sext = {{11{imm_j[20]}}, imm_j[20:0]};

  // opcodes - see section 19 of RiscV spec
  localparam bit [`OPCODE_SIZE] OpLoad = 7'b00_000_11;
  localparam bit [`OPCODE_SIZE] OpStore = 7'b01_000_11;
  localparam bit [`OPCODE_SIZE] OpBranch = 7'b11_000_11;
  localparam bit [`OPCODE_SIZE] OpJalr = 7'b11_001_11;
  localparam bit [`OPCODE_SIZE] OpMiscMem = 7'b00_011_11;
  localparam bit [`OPCODE_SIZE] OpJal = 7'b11_011_11;

  localparam bit [`OPCODE_SIZE] OpRegImm = 7'b00_100_11;
  localparam bit [`OPCODE_SIZE] OpRegReg = 7'b01_100_11;
  localparam bit [`OPCODE_SIZE] OpEnviron = 7'b11_100_11;

  localparam bit [`OPCODE_SIZE] OpAuipc = 7'b00_101_11;
  localparam bit [`OPCODE_SIZE] OpLui = 7'b01_101_11;

  wire insn_lui = insn_opcode == OpLui;
  wire insn_auipc = insn_opcode == OpAuipc;
  wire insn_jal = insn_opcode == OpJal;
  wire insn_jalr = insn_opcode == OpJalr;

  wire insn_beq = insn_opcode == OpBranch && insn_from_imem[14:12] == 3'b000;
  wire insn_bne = insn_opcode == OpBranch && insn_from_imem[14:12] == 3'b001;
  wire insn_blt = insn_opcode == OpBranch && insn_from_imem[14:12] == 3'b100;
  wire insn_bge = insn_opcode == OpBranch && insn_from_imem[14:12] == 3'b101;
  wire insn_bltu = insn_opcode == OpBranch && insn_from_imem[14:12] == 3'b110;
  wire insn_bgeu = insn_opcode == OpBranch && insn_from_imem[14:12] == 3'b111;

  wire insn_lb = insn_opcode == OpLoad && insn_from_imem[14:12] == 3'b000;
  wire insn_lh = insn_opcode == OpLoad && insn_from_imem[14:12] == 3'b001;
  wire insn_lw = insn_opcode == OpLoad && insn_from_imem[14:12] == 3'b010;
  wire insn_lbu = insn_opcode == OpLoad && insn_from_imem[14:12] == 3'b100;
  wire insn_lhu = insn_opcode == OpLoad && insn_from_imem[14:12] == 3'b101;

  wire insn_sb = insn_opcode == OpStore && insn_from_imem[14:12] == 3'b000;
  wire insn_sh = insn_opcode == OpStore && insn_from_imem[14:12] == 3'b001;
  wire insn_sw = insn_opcode == OpStore && insn_from_imem[14:12] == 3'b010;

  wire insn_addi = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b000;
  wire insn_slti = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b010;
  wire insn_sltiu = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b011;
  wire insn_xori = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b100;
  wire insn_ori = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b110;
  wire insn_andi = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b111;

  wire insn_slli = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b001 && insn_from_imem[31:25] == 7'd0;
  wire insn_srli = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b101 && insn_from_imem[31:25] == 7'd0;
  wire insn_srai = insn_opcode == OpRegImm && insn_from_imem[14:12] == 3'b101 && insn_from_imem[31:25] == 7'b0100000;

  wire insn_add = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b000 && insn_from_imem[31:25] == 7'd0;
  wire insn_sub  = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b000 && insn_from_imem[31:25] == 7'b0100000;
  wire insn_sll = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b001 && insn_from_imem[31:25] == 7'd0;
  wire insn_slt = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b010 && insn_from_imem[31:25] == 7'd0;
  wire insn_sltu = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b011 && insn_from_imem[31:25] == 7'd0;
  wire insn_xor = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b100 && insn_from_imem[31:25] == 7'd0;
  wire insn_srl = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b101 && insn_from_imem[31:25] == 7'd0;
  wire insn_sra  = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b101 && insn_from_imem[31:25] == 7'b0100000;
  wire insn_or = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b110 && insn_from_imem[31:25] == 7'd0;
  wire insn_and = insn_opcode == OpRegReg && insn_from_imem[14:12] == 3'b111 && insn_from_imem[31:25] == 7'd0;

  wire insn_mul    = insn_opcode == OpRegReg && insn_from_imem[31:25] == 7'd1 && insn_from_imem[14:12] == 3'b000;
  wire insn_mulh   = insn_opcode == OpRegReg && insn_from_imem[31:25] == 7'd1 && insn_from_imem[14:12] == 3'b001;
  wire insn_mulhsu = insn_opcode == OpRegReg && insn_from_imem[31:25] == 7'd1 && insn_from_imem[14:12] == 3'b010;
  wire insn_mulhu  = insn_opcode == OpRegReg && insn_from_imem[31:25] == 7'd1 && insn_from_imem[14:12] == 3'b011;
  wire insn_div    = insn_opcode == OpRegReg && insn_from_imem[31:25] == 7'd1 && insn_from_imem[14:12] == 3'b100;
  wire insn_divu   = insn_opcode == OpRegReg && insn_from_imem[31:25] == 7'd1 && insn_from_imem[14:12] == 3'b101;
  wire insn_rem    = insn_opcode == OpRegReg && insn_from_imem[31:25] == 7'd1 && insn_from_imem[14:12] == 3'b110;
  wire insn_remu   = insn_opcode == OpRegReg && insn_from_imem[31:25] == 7'd1 && insn_from_imem[14:12] == 3'b111;

  wire insn_ecall = insn_opcode == OpEnviron && insn_from_imem[31:7] == 25'd0;
  wire insn_fence = insn_opcode == OpMiscMem;

  // synthesis translate_off
  // this code is only for simulation, not synthesis
  `include "RvDisassembler.sv"
  string disasm_string;
  always_comb begin
    disasm_string = rv_disasm(insn_from_imem);
  end
  // HACK: get disasm_string to appear in GtkWave, which can apparently show only wire/logic...
  wire [(8*32)-1:0] disasm_wire;
  genvar i;
  for (i = 0; i < 32; i = i + 1) begin : gen_disasm
    assign disasm_wire[(((i+1))*8)-1:((i)*8)] = disasm_string[31-i];
  end
  // synthesis translate_on

  // program counter
  logic [`REG_SIZE] pcNext, pcCurrent;
  always @(posedge clk) begin
    if (rst) begin
      pcCurrent <= 32'd0;
    end else begin
      pcCurrent <= pcNext;
    end
  end
  assign pc_to_imem = pcCurrent;

  // cycle/insn_from_imem counters
  logic [`REG_SIZE] cycles_current, num_insns_current;
  always @(posedge clk) begin
    if (rst) begin
      cycles_current <= 0;
      num_insns_current <= 0;
    end else begin
      cycles_current <= cycles_current + 1;
      if (!rst) begin
        num_insns_current <= num_insns_current + 1;
      end
    end
  end

  logic illegal_insn;
  logic we; 
  logic [4:0]rs1;
  logic [4:0]rs2;
  logic [4:0]rd;
  logic [31:0]rs2_data;
  logic [31:0]rs1_data;
  logic [31:0]rd_data;
  logic [31:0]imm;
  logic [31:0] signextended;
  logic [6:0] func7;
  logic [12:0] offset;
  logic [12:0] offsetshift;
  logic [20:0] targ20;
  RegFile rf(.rd(rd), .rd_data(rd_data), .rs1(rs1), .rs1_data(rs1_data), .rs2(rs2), .rs2_data(rs2_data), .clk(clk), .we(we), .rst(rst));

  logic [31:0]inputone; 
  logic [31:0]inputtwo;
  logic [2:0] fun3;
  logic [6:0] fun7;
  logic [6:0] opcode;
  logic [31:0] aluresult;
  logic signeddivflag;

  ALU al(.inputone(inputone), .inputtwo(inputtwo), .opcode(opcode), .fun3(fun3), .fun7(fun7), .signeddivflag(signeddivflag), .aluresult(aluresult));


  always_comb begin
    illegal_insn = 1'b0;
    halt = 0;
    we = 1'b0;
    case (insn_opcode)
      OpLui: begin
        opcode = insn_opcode;
        we = 1'b1;
        rd = insn_from_imem[11:7];
        rd_data = {insn_from_imem[31:12], 12'b0};
        pcNext = pcCurrent + 32'd4;
      end

      OpAuipc: begin
        opcode = insn_opcode;
        we = 1'b1;
        rd = insn_from_imem[11:7];
        rd_data = pcCurrent + {insn_from_imem[31:12], 12'b0};
        pcNext = pcCurrent + 32'd4;
      end

      OpRegImm: begin
        opcode = insn_opcode;
        we = 1'b1;
        rs1 = insn_from_imem[19:15];
        rd = insn_from_imem[11:7];
        fun3 =insn_from_imem[14:12];

        case(insn_from_imem[14:12]) 
        3'b000: begin
          imm[11:0] = insn_from_imem[31:20];
          signextended = {{20{imm[11]}},imm[11:0]};
          inputone = rs1_data;
          inputtwo = signextended;
          rd_data = aluresult;
        end
        3'b010: begin
          imm[11:0] = insn_from_imem[31:20];
          signextended = {{20{imm[11]}},imm[11:0]};
          inputone = rs1_data;
          inputtwo = signextended;
          rd_data = aluresult;
        end

        3'b011: begin 
          imm[11:0] = insn_from_imem[31:20];
          signextended = {{20{imm[11]}},imm[11:0]};
          inputone = rs1_data;
          inputtwo = signextended;
          rd_data = aluresult;
        end

        3'b100: begin 
          imm[11:0] = insn_from_imem[31:20];
          signextended = {{20{imm[11]}},imm[11:0]};
          inputone = rs1_data;
          inputtwo = signextended;
          rd_data = aluresult;
        end

        3'b110: begin 
          imm[11:0] = insn_from_imem[31:20];
          signextended = {{20{imm[11]}},imm[11:0]};
          inputone = rs1_data;
          inputtwo = signextended;
          rd_data = aluresult;
        end

        3'b111: begin 
          imm[11:0] = insn_from_imem[31:20];
          signextended = {{20{imm[11]}},imm[11:0]};
          inputone = rs1_data;
          inputtwo = signextended;
          rd_data = aluresult;
        end

        3'b001: begin 
          rd_data = rs1_data << insn_from_imem[24:20];
        end

        3'b101: begin 
          if(insn_from_imem[31:25]==7'd0) begin
            rd_data = rs1_data >> insn_from_imem[24:20];
          end
          if(insn_from_imem[31:25]==7'd32) begin
            rd_data = $signed(rs1_data) >>> insn_from_imem[24:20];
          end
        end        
        default: begin
        end
        endcase
        pcNext = pcCurrent + 32'd4;

      end

      OpRegReg: begin
      opcode = insn_opcode;
      we = 1'b1;
      rs1 = insn_from_imem[19:15];
      rs2 = insn_from_imem[24:20];
      rd = insn_from_imem[11:7];
      inputone = rs1_data;
      fun7 = insn_from_imem[31:25];        
      fun3 =insn_from_imem[14:12];
       case(insn_from_imem[14:12])
       3'b000: begin
        if(fun7==7'd0) begin
          inputtwo = rs2_data;
        end
        if(fun7==7'd1) begin
          inputtwo = rs2_data;
        end
        if(fun7==7'd32) begin
          inputtwo = ~rs2_data;
        end
        rd_data = aluresult;
       end

       3'b100: begin
        if (fun7 == 7'd1) begin
          inputone = rs1_data[31] == 0 ? rs1_data : ~(rs1_data) + 1;
          inputtwo = rs2_data[31] == 0 ? rs2_data : ~(rs2_data) + 1;
          signeddivflag = rs1_data[31] != rs2_data[31];
        end else begin
          inputone = rs1_data;
          inputtwo = rs2_data;
        end
        rd_data = aluresult;
       end

       3'b110: begin
        if (fun7 == 7'd1) begin
          inputone = rs1_data[31] == 0 ? rs1_data : ~(rs1_data) + 1;
          inputtwo = rs2_data[31] == 0 ? rs2_data : ~(rs2_data) + 1;
          signeddivflag = rs1_data[31] == 1'b1;
        end else begin
          inputone = rs1_data;
          inputtwo = rs2_data;
        end
        rd_data = aluresult;
       end
      
      default: begin 
        inputone = rs1_data;
        inputtwo = rs2_data;
        rd_data = aluresult;
      end
      endcase
      pcNext = pcCurrent + 32'd4;
      end

      OpEnviron: 
        begin
          halt = 1;
          pcNext = pcCurrent + 32'd4;
        end
      
      OpBranch:
      begin
      offset[12] = insn_from_imem[31];
      offset[10:5] = insn_from_imem[30:25];
      offset[4:1] = insn_from_imem[11:8];
      offset[11] = insn_from_imem[7];
      offset[0] = 0;
      offsetshift = offset;
      imm = {{19{offsetshift[12]}}, offsetshift[12:0]};
      rs1 = insn_from_imem[19:15];
      rs2 = insn_from_imem[24:20];
        
        case(insn_from_imem[14:12])
       3'b000: begin
        if(rs1_data == rs2_data) begin
          inputone = pcCurrent;
          inputtwo = imm;
          fun3 = 3'b0;
          opcode = OpRegImm;
          pcNext = aluresult;
        end else begin
          pcNext = pcCurrent + 32'd4;
        end
       end

       3'b001: begin
        if(rs1_data != rs2_data) begin
          inputone = pcCurrent;
          inputtwo = imm;
          fun3 = 3'b0;
          opcode = OpRegImm;
          pcNext = aluresult;
        end else begin
          pcNext = pcCurrent + 32'd4;
        end
       end

        3'b100: begin
        if($signed(rs1_data) < $signed(rs2_data)) begin
          inputone = pcCurrent;
          inputtwo = imm;
          fun3 = 3'b0;
          opcode = OpRegImm;
          pcNext = aluresult;
        end else begin
          pcNext = pcCurrent + 32'd4;
        end
       end

        3'b101: begin
        if($signed(rs1_data) >= $signed(rs2_data)) begin
          inputone = pcCurrent;
          inputtwo = imm;
          fun3 = 3'b0;
          opcode = OpRegImm;
          pcNext = aluresult;
        end else begin
          pcNext = pcCurrent + 32'd4;
        end
       end

        3'b110: begin
        if(rs1_data < rs2_data) begin
          inputone = pcCurrent;
          inputtwo = imm;
          fun3 = 3'b0;
          opcode = OpRegImm;
          pcNext = aluresult;
        end else begin
          pcNext = pcCurrent + 32'd4;
        end
       end

       3'b111: begin
        if(rs1_data >= rs2_data) begin
          inputone = pcCurrent;
          inputtwo = imm;
          fun3 = 3'b0;
          opcode = OpRegImm;
          pcNext = aluresult;
        end else begin
          pcNext = pcCurrent + 32'd4;
        end
       end
        default: begin end
        endcase
       end

       OpJal: begin
          targ20[20] = insn_from_imem[31];
          targ20[10:1] = insn_from_imem[30:21];
          targ20[11] = insn_from_imem[20];
          targ20[19:12] = insn_from_imem[19:12];
          targ20[0] = 0;
          opcode = OpJal;
          inputone = pcCurrent;
          inputtwo = {{11{targ20[20]}}, targ20[20:0]};
          pcNext = aluresult;
          we = 1'b1;
          rd = insn_from_imem[11:7];
          rd_data = pcCurrent + 32'd4;
       end

       OpJalr: begin
          we = 1'b1;
          rd = insn_from_imem[11:7];
          rd_data = pcCurrent + 32'd4;
          rs1 = insn_from_imem[19:15];
          pcNext = ((rs1_data + {{20{insn_from_imem[31]}}, insn_from_imem[31:20]}) & ~32'b1);
       end

       OpLoad: begin
        opcode = insn_opcode;
        fun3 = insn_from_imem[14:12];
        we = 1'b1;
        rd = insn_from_imem[11:7];
        rs1 = insn_from_imem[19:15];
        pcNext = pcCurrent + 32'd4;
        store_we_to_dmem = 4'b0;
        addr_to_dmem = (rs1_data + {{20{insn_from_imem[31]}}, insn_from_imem[31:20]}) & {{30{1'b1}},{2{1'b0}}};
        inputone = load_data_from_dmem;
        inputtwo = ((rs1_data + {{20{insn_from_imem[31]}}, insn_from_imem[31:20]}) << 3) & {{27{1'b0}}, {2{1'b1}} , {3{1'b0}}};
        rd_data = aluresult;
       end

       OpStore: begin
        opcode = insn_opcode;
        fun3 = insn_from_imem[14:12];
        we = 1'b0;
        pcNext = pcCurrent + 32'd4;
        rs1 = insn_from_imem[19:15];
        rs2 = insn_from_imem[24:20];
        imm = rs1_data + {{20{insn_from_imem[31]}}, insn_from_imem[31:25], insn_from_imem[11:7]};
        
        case (fun3)
          3'b000: begin
            store_we_to_dmem = 4'b1 << imm[1:0];
            addr_to_dmem = imm & {{30{1'b1}},{2{1'b0}}};
            store_data_to_dmem = rs2_data << {imm[1:0], 3'b0};
          end
          3'b001: begin
            store_we_to_dmem = 4'b11 << imm[1:0];
            addr_to_dmem = imm & {{30{1'b1}},{2{1'b0}}};
            store_data_to_dmem = rs2_data << {imm[1:0], 3'b0};
          end
          3'b010: begin
            store_we_to_dmem = 4'b1111;
            addr_to_dmem = imm & {{30{1'b1}},{2{1'b0}}};
            store_data_to_dmem = rs2_data << {imm[1:0], 3'b0};
          end
          default: begin end

        endcase
       end

      default: begin
        illegal_insn = 1'b1;
        pcNext = pcCurrent + 32'd4;
      end

    endcase
  end

endmodule

module ALU (
  input logic [31:0]inputone,
  input logic [31:0]inputtwo,
  input logic [2:0]fun3,
  input logic [6:0]opcode,
  input logic [6:0]fun7,
  input logic signeddivflag,
  output logic [31:0] aluresult
);
logic [31:0] claoutput;
logic [31:0] quotient;
logic [31:0] remainder;
logic cin;
cla cla(.a(inputone), .b(inputtwo), .cin(cin), .sum(claoutput));
divider_unsigned div(.i_dividend(inputone), .i_divisor(inputtwo), .o_quotient(quotient), .o_remainder(remainder));

logic [63:0] mulresult;
logic [31:0] memaddress;

always_comb begin
case(opcode)
7'b00_100_11: begin
  case(fun3)
  3'b000: begin 
    cin=0;
    aluresult = claoutput;
  end

  3'b010: begin 
    if($signed(inputone) < $signed(inputtwo)) begin
      aluresult = 1;
    end else begin
      aluresult = 0;
    end
  end

  3'b011: begin 
    if(inputone < inputtwo) begin
      aluresult = 1;
    end else begin
      aluresult = 0;
    end
  end

  3'b100: begin 
    aluresult = inputone ^ inputtwo;
  end

  3'b110: begin 
    aluresult = inputone | inputtwo;
  end

  3'b111: begin 
    aluresult = inputone & inputtwo;
  end

  default: begin end
  endcase
end

7'b11_011_11: begin
  cin = 0;
  aluresult = claoutput;
end

7'b00_000_11: begin
  case(fun3)
    3'b000: begin
      memaddress = (inputone >> inputtwo[4:0]);
      aluresult = {{24{memaddress[7]}}, memaddress[7:0]};
    end
    3'b001: begin
      memaddress = (inputone >> inputtwo[4:0]);
      aluresult = {{16{memaddress[15]}}, memaddress[15:0]};
    end
    3'b010: begin
      memaddress = (inputone >> inputtwo[4:0]);
      aluresult = memaddress;
    end
    3'b100: begin
      memaddress = (inputone >> inputtwo[4:0]);
      aluresult = {24'b0, memaddress[7:0]};
    end
    3'b101: begin
      memaddress = (inputone >> inputtwo[4:0]);
      aluresult = {16'b0, memaddress[15:0]};
    end
    default: begin end
  endcase
  
end

7'b01_100_11: begin
  case(fun3)
  3'b000: begin 
    case(fun7)
    7'd0: begin 
      cin = 0;
      aluresult = claoutput;
    end
    7'd1: begin
      mulresult = inputone * inputtwo;
      aluresult = mulresult[31:0];
    end
    7'd32: begin 
      cin = 1;
      aluresult = claoutput;
    end
    default: begin 
      aluresult = claoutput;
    end
    endcase
  end

  3'b001: begin
    case (fun7)
      7'd0: begin
        aluresult = inputone << inputtwo[4:0];
      end
      7'd1: begin
        mulresult = $signed(inputone) * $signed(inputtwo);
        aluresult = mulresult[63:32];
      end
      default: begin
        aluresult = claoutput;
      end
    endcase
  end

  3'b010: begin 
    case (fun7)
      7'd0: begin
        if($signed(inputone) < $signed(inputtwo)) begin
          aluresult = 1;
        end else begin
          aluresult = 0;
        end
      end
      7'd1: begin
        mulresult = {{32{inputone[31]}}, inputone[31:0]} * {32'b0, inputtwo[31:0]};
        aluresult = mulresult[63:32];
      end
      default: begin
        aluresult = claoutput;
      end
    endcase
  end

  3'b011: begin 
    case (fun7)
      7'd0: begin
        if(inputone < inputtwo) begin
          aluresult = 1;
        end else begin
          aluresult = 0;
        end
      end
      7'd1: begin
        mulresult = inputone * inputtwo;
        aluresult = mulresult[63:32];
      end
      default: begin
        aluresult = claoutput;
      end
    endcase
  end

  3'b100: begin 
    case (fun7)
      7'd0: begin
        aluresult = inputone ^ inputtwo;
      end
      7'd1: begin
        aluresult = inputtwo == 32'b0 ? ({32{1'b1}}) : (signeddivflag ? ~(quotient) + 1 : quotient);
      end
      default: begin
        aluresult = claoutput;
      end
    endcase
    
  end

  3'b101: begin 
          if(fun7==7'd0) begin
            aluresult = inputone >> inputtwo[4:0];
          end
          if(fun7==7'd1) begin
            aluresult = quotient;
          end
          if(fun7==7'd32) begin
            aluresult = $signed(inputone) >>> inputtwo[4:0];
          end
  end

  3'b110: begin 
    case (fun7)
      7'd0: begin
        aluresult = inputone | inputtwo;
      end
      7'd1: begin
        aluresult = inputtwo == 32'b0 ? (inputone == 32'b0 ? 32'b0 : (signeddivflag ? {1'b1, 31'b0} : 32'b1)) : (signeddivflag ? ~(remainder) + 1 : remainder);
      end
      default: begin
        aluresult = claoutput;
      end
    endcase
  end

  3'b111: begin 
    if(fun7==7'd0) begin
      aluresult = inputone & inputtwo;
    end
    if(fun7==7'd1) begin
      aluresult = remainder;
    end
  end

  default: begin end
  endcase
end


default: begin end
endcase
end
endmodule

/* A memory module that supports 1-cycle reads and writes, with one read-only port
 * and one read+write port.
 */
module MemorySingleCycle #(
    parameter int NUM_WORDS = 512
) (
    // rst for both imem and dmem
    input wire rst,

    // clock for both imem and dmem. See RiscvProcessor for clock details.
    input wire clock_mem,

    // must always be aligned to a 4B boundary
    input wire [`REG_SIZE] pc_to_imem,

    // the value at memory location pc_to_imem
    output logic [`REG_SIZE] insn_from_imem,

    // must always be aligned to a 4B boundary
    input wire [`REG_SIZE] addr_to_dmem,

    // the value at memory location addr_to_dmem
    output logic [`REG_SIZE] load_data_from_dmem,

    // the value to be written to addr_to_dmem, controlled by store_we_to_dmem
    input wire [`REG_SIZE] store_data_to_dmem,

    // Each bit determines whether to write the corresponding byte of store_data_to_dmem to memory location addr_to_dmem.
    // E.g., 4'b1111 will write 4 bytes. 4'b0001 will write only the least-significant byte.
    input wire [3:0] store_we_to_dmem
);

  // memory is arranged as an array of 4B words
  logic [`REG_SIZE] mem[NUM_WORDS];

  initial begin
    $readmemh("mem_initial_contents.hex", mem, 0);
  end

  always_comb begin
    // memory addresses should always be 4B-aligned
    assert (pc_to_imem[1:0] == 2'b00);
    assert (addr_to_dmem[1:0] == 2'b00);
  end

  localparam int AddrMsb = $clog2(NUM_WORDS) + 1;
  localparam int AddrLsb = 2;

  always @(posedge clock_mem) begin
    if (rst) begin
    end else begin
      insn_from_imem <= mem[{pc_to_imem[AddrMsb:AddrLsb]}];
    end
  end

  always @(negedge clock_mem) begin
    if (rst) begin
    end else begin
      if (store_we_to_dmem[0]) begin
        mem[addr_to_dmem[AddrMsb:AddrLsb]][7:0] <= store_data_to_dmem[7:0];
      end
      if (store_we_to_dmem[1]) begin
        mem[addr_to_dmem[AddrMsb:AddrLsb]][15:8] <= store_data_to_dmem[15:8];
      end
      if (store_we_to_dmem[2]) begin
        mem[addr_to_dmem[AddrMsb:AddrLsb]][23:16] <= store_data_to_dmem[23:16];
      end
      if (store_we_to_dmem[3]) begin
        mem[addr_to_dmem[AddrMsb:AddrLsb]][31:24] <= store_data_to_dmem[31:24];
      end
      // dmem is "read-first": read returns value before the write
      load_data_from_dmem <= mem[{addr_to_dmem[AddrMsb:AddrLsb]}];
    end
  end
endmodule

/*
This shows the relationship between clock_proc and clock_mem. The clock_mem is
phase-shifted 90° from clock_proc. You could think of one proc cycle being
broken down into 3 parts. During part 1 (which starts @posedge clock_proc)
the current PC is sent to the imem. In part 2 (starting @posedge clock_mem) we
read from imem. In part 3 (starting @negedge clock_mem) we read/write memory and
prepare register/PC updates, which occur at @posedge clock_proc.

        ____
 proc: |    |______
           ____
 mem:  ___|    |___
*/
module RiscvProcessor (
    input  wire  clock_proc,
    input  wire  clock_mem,
    input  wire  rst,
    output logic halt
);

  wire [`REG_SIZE] pc_to_imem, insn_from_imem, mem_data_addr, mem_data_loaded_value, mem_data_to_write;
  wire [3:0] mem_data_we;

  MemorySingleCycle #(
      .NUM_WORDS(8192)
  ) mem (
      .rst      (rst),
      .clock_mem (clock_mem),
      // imem is read-only
      .pc_to_imem(pc_to_imem),
      .insn_from_imem(insn_from_imem),
      // dmem is read-write
      .addr_to_dmem(mem_data_addr),
      .load_data_from_dmem(mem_data_loaded_value),
      .store_data_to_dmem (mem_data_to_write),
      .store_we_to_dmem  (mem_data_we)
  );

  DatapathSingleCycle datapath (
      .clk(clock_proc),
      .rst(rst),
      .pc_to_imem(pc_to_imem),
      .insn_from_imem(insn_from_imem),
      .addr_to_dmem(mem_data_addr),
      .store_data_to_dmem(mem_data_to_write),
      .store_we_to_dmem(mem_data_we),
      .load_data_from_dmem(mem_data_loaded_value),
      .halt(halt)
  );

endmodule
